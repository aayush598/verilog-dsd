module NOT_gate (A,Y);
	input A;
	output Y;
	assign Y = ~A;
endmodule