module XOR_gate(
	input wire A,
	input wire B,
	output reg Y);

	assign Y = A^B;

endmodule